module register_file (s, enable, load, reset, clock, selectA, selectB, MA, MB);
input [0:4] s;
input enable, load, reset, clock;
input [0:4] selectA;
input [0:4] selectB;
output reg [0:31] MA, MB;
endmodule

module decoder(s,enable,I);
input [0:4] s;
input enable;
output reg [0:31] I;

always @(s or enable)
begin
	if (enable == 0)
		I = 32'b00000000000000000000000000000000;
		
	else
		case(s)
			5'b00000: I = 32'b00000000000000000000000000000001;
			5'b00001: I = 32'b00000000000000000000000000000010;
			5'b00010: I = 32'b00000000000000000000000000000100;
			5'b00011: I = 32'b00000000000000000000000000001000;
			5'b00100: I = 32'b00000000000000000000000000010000;
			5'b00101: I = 32'b00000000000000000000000000100000;
			5'b00110: I = 32'b00000000000000000000000001000000;
			5'b00111: I = 32'b00000000000000000000000010000000;
			5'b01000: I = 32'b00000000000000000000000100000000;
			5'b01001: I = 32'b00000000000000000000001000000000;
			5'b01010: I = 32'b00000000000000000000010000000000;
			5'b01011: I = 32'b00000000000000000000100000000000;
			5'b01100: I = 32'b00000000000000000001000000000000;
			5'b01101: I = 32'b00000000000000000010000000000000;
			5'b01110: I = 32'b00000000000000000100000000000000;
			5'b01111: I = 32'b00000000000000001000000000000000;
			5'b10000: I = 32'b00000000000000010000000000000000;
			5'b10001: I = 32'b00000000000000100000000000000000;
			5'b10010: I = 32'b00000000000001000000000000000000; 
			5'b10011: I = 32'b00000000000010000000000000000000;
			5'b10100: I = 32'b00000000000100000000000000000000;
			5'b10101: I = 32'b00000000001000000000000000000000;
			5'b10110: I = 32'b00000000010000000000000000000000;
			5'b10111: I = 32'b00000000100000000000000000000000;
			5'b11000: I = 32'b00000001000000000000000000000000;
			5'b11001: I = 32'b00000010000000000000000000000000;
			5'b11010: I = 32'b00000100000000000000000000000000;
			5'b11011: I = 32'b00001000000000000000000000000000;
			5'b11100: I = 32'b00010000000000000000000000000000;
			5'b11101: I = 32'b00100000000000000000000000000000;
			5'b11110: I = 32'b01000000000000000000000000000000;
			5'b11111: I = 32'b10000000000000000000000000000000;
		default I = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
		endcase
	end
endmodule

module register(I,clock,reset,load,O);
input [0:31] I;
input load;
input clock;
input reset;
output reg [0:31] O;

always @(posedge clock)
begin
	if (reset == 1)
		O <= 0;
	else
	if (load == 1)
		O <= I;
		end
endmodule

module muxA(O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31,selectA,MA);

parameter N=32;
input [N-1:0] O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31;
input [0:4] selectA;
output reg [N-1:0] MA;


always @(O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31 or selectA)
begin
	case(selectA)
		5'b00000: MA = O0;
		5'b00001: MA = O1;
		5'b00010: MA = O2;
		5'b00011: MA = O3;
		5'b00100: MA = O4;
		5'b00101: MA = O5;
		5'b00110: MA = O6;
		5'b00111: MA = O7;
		5'b01000: MA = O8;
		5'b01001: MA = O9;
		5'b01010: MA = O10;
		5'b01011: MA = O11;
		5'b01100: MA = O12;
		5'b01101: MA = O13;
		5'b01110: MA = O14;
		5'b01111: MA = O15;
		5'b10000: MA = O16;
		5'b10001: MA = O17;
		5'b10010: MA = O18;
		5'b10011: MA = O19;
		5'b10100: MA = O20;
		5'b10101: MA = O21;
		5'b10110: MA = O22;
		5'b10111: MA = O23;
		5'b11000: MA = O24;
		5'b11001: MA = O25;
		5'b11010: MA = O26;
		5'b11011: MA = O27;
		5'b11100: MA = O28;
		5'b11101: MA = O29;
		5'b11110: MA = O30;
		5'b11111: MA = O31;
		default MA = 1'bx;
	endcase
	end
endmodule

module muxB(O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31,selectB,MB);

parameter N=32;
input [N-1:0] O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31;
input [0:4] selectB;
output reg [N-1:0] MB;


always @(O0,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31 or selectB)
begin
	case(selectB)
		5'b00000: MB = O0;
		5'b00001: MB = O1;
		5'b00010: MB = O2;
		5'b00011: MB = O3;
		5'b00100: MB = O4;
		5'b00101: MB = O5;
		5'b00110: MB = O6;
		5'b00111: MB = O7;
		5'b01000: MB = O8;
		5'b01001: MB = O9;
		5'b01010: MB = O10;
		5'b01011: MB = O11;
		5'b01100: MB = O12;
		5'b01101: MB = O13;
		5'b01110: MB = O14;
		5'b01111: MB = O15;
		5'b10000: MB = O16;
		5'b10001: MB = O17;
		5'b10010: MB = O18;
		5'b10011: MB = O19;
		5'b10100: MB = O20;
		5'b10101: MB = O21;
		5'b10110: MB = O22;
		5'b10111: MB = O23;
		5'b11000: MB = O24;
		5'b11001: MB = O25;
		5'b11010: MB = O26;
		5'b11011: MB = O27;
		5'b11100: MB = O28;
		5'b11101: MB = O29;
		5'b11110: MB = O30;
		5'b11111: MB = O31;
		default MB = 1'bx;
	endcase
	end
endmodule

